-- Memoria de instruciones 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

entity mem_inst is
generic (n: natural:=8); -- n�mero de bits de direcci�n
port (
-- direcci�n de lectura/escritura
dir : in std_logic_vector(n-1 downto 0); 
dout : out std_logic_vector(31 downto 0));
end mem_inst;

architecture compor of mem_inst is
type rom_type is array (0 to 2**n - 1) of std_logic_vector (7 downto 0);
-- la se�al RAM puede inicializarse asign�ndole valores.
signal RAM: rom_type:= (X"00", "00000100", -- 0
"00011000", "00100010", -- Sub $3, $0, $4
"10101100", "00000100", -- 4	
"00000000", "00001000", -- Sw $4, 8($0)
"00000000", "00000000", -- 8
"00000000", "00000000", -- nop 
"00100000", "01100001", -- 12
"00000000", "00010111", -- addi $1, $3, 23
"00101000", "01101000", -- 16
"11111111", "11111110", -- slti $8, $3, -2 
"00000000", "00000000", -- 20
"00000000", "00000000", -- nop 
"00000000", "00100011", -- 24
"00010000", "00100100", -- And $2, $1, $3 
"00000001", "00000011", -- 28	
"00101000", "00100111", -- Nor $5, $8, $3
"10001100", "00000110", -- 32	
"00000000", "00010100", -- Lw $6, 20($0) 
"00001100", "00000000", -- 36	
"00000000", "01100100", -- Jal rutina : dir=100

--Hecho por nosotros
"00000000", "00000000", -- 40
"00000000", "00000000", -- nop 
"10101100", "00000010", -- 44
"00000000", "00001100", -- Sw $2, 12($0)
"10101100", "00001000", -- 48
"00000000", "00001000", -- Sw $8, 8($0)
"10101100", "00000101", -- 52
"00000000", "00000100", -- Sw $5, 4($0)
"10001100", "00001001", -- 56
"00000000", "00001100", -- Lw $9, 12($0)
"00000000", "00000000", -- 60
"00000000", "00000000", -- nop 
"00000000", "00000000", -- 64
"00000000", "00000000", -- nop 
"00000001", "00101000",	-- 68
"00001000", "00100010", -- Sub $1, $9, $8
"00010100", "00000011", -- 72 = fin
"11111111", "11111111", -- Bne $0, $3, -1
"00000000", "00000000", -- 76
"00000000", "00000000", -- nop 

"00000000", "00000000", -- 80
"00000000", "00000000", -- nop 
"00000000", "00000000", -- 84
"00000000", "00000000", -- nop 
"00000000", "00000000", -- 88
"00000000", "00000000", -- nop 
"00000000", "00000000", -- 92
"00000000", "00000000", -- nop 
"00000000", "00000000", -- 96
"00000000", "00000000", -- nop 

"00000000", "00100001", -- 100 = rutina
"00011000", "00100110", -- xor $3,$1,$1
"00110100", "00000010", -- 104
"00000000", "00000000", -- Ori $2, $0, 0
"00000000", "00000000", -- 108
"00000000", "00000000", -- nop
"00000000", "01100110", -- 112 = bucle
"00001000", "00101010", -- slt $1, $3, $6
"00000000", "00000000", -- 116
"00000000", "00000000", -- nop
"00000000", "00000000", -- 120
"00000000", "00000000", -- nop
"00010000", "00100000", -- 124
--fin de lo nuestro


"00000000", "00000110", -- Beq $1, $0, ret
"00000000", "00000000", -- 128
"00000000", "00000000", -- nop 
"10001100", "10000101", -- 132	
"00000000", "00000000", -- Lw $5, 0($4) 
"00100000", "01100011", -- 136
"00000000", "00000001", -- Addi $3, $3, 1
"00100000", "10000100", -- 140
"00000000", "00000100", -- Addi $4, $4, 4
"00001000", "00000000", -- 144
"00000000", "01110000", -- J bucle = 112
"00000000", "01000101", -- 148
"00010000", "00100000", -- Add $2, $2, $5 (hueco relleno)
"00000001", "11100000", -- 152 = ret
"00000000", "00001000", -- jr $15 
"00000000", "00000000", -- 156
"00000000", "00000000", -- nop 
others => X"00");

signal MSB, M3B,m2b, LSB: std_logic_vector(7 downto 0);

Begin

-- proceso de lectura as�ncrona	
MSB <= RAM(conv_integer(dir));
M2b <= RAM(conv_integer(dir + 1));
m3b <= RAM(conv_integer(dir + 2));
LSB <= RAM(conv_integer(dir + 3));
dout <= MSB & M2b & m3b & LSB;
end compor;